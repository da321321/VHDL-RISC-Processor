-------------------------------------------------------------------------------
-- ubus
-- by fcampi@sfu.ca Feb 2014
--
-- Local Bus for the internal data bus
-- of the Qrisc processor up island
-------------------------------------------------------------------------------

-- There is an interesting challenge in this design, that is how to handle
-- ready signals coming from the slaves in case slaves have a response time
-- higher than 1 cycle, for example FIFOs that may be empty or full.
-- The bus is based on 2 main cycles: the addressing cycle C1, and the reading
-- cycle C2 separated by a clock.
-- 
-- Note: 
-- NREADY is generated BY A SLAVE to A BUS, when it is not able to respond to the bus request
-- (example, a multicyle memory saying "I am not ready yet")
-- BUSY  is generated BY A MASTER, when it needs an extension of the current
-- bus cyle (Example, the master is stalled and is in no condition to read incoming data)

-- NREADY when fed to a master can be due to many different configurations:
-- -- a) Master is requiring the bus but another master is having it
   -- b) The slave addressed by the master needs an extension during the addressing
   -- c) The Master in charge of the previous bus run needs an extension during reading


library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

  entity ubus is
    generic(signal_active : std_logic := '0';
            addr_size : positive := 32; size : positive := 32; -- need to edit it to 16 bits
            s1_start  : Std_logic_vector := X"40001000";
            s1_end    : Std_logic_vector := X"40002000";
            s2_start  : Std_logic_vector := X"50000000";
            s2_end    : Std_logic_vector := X"f0000000";
            s3_start  : Std_logic_vector := X"00000000";
            s3_end    : Std_logic_vector := X"00000000";
            s4_start  : Std_logic_vector := X"00000000";
            s4_end    : Std_logic_vector := X"00000000" );
      
    port ( clk,reset           : in Std_logic;
           -- M1 port
           M1_BUSY,M1_MR,M1_MW : in   Std_logic;
           M1_NREADY           : out  Std_logic;
           M1_ADDRBUS          : in   Std_logic_vector(addr_size-1 downto 0);
           M1_RDATABUS         : out  Std_logic_vector(size-1 downto 0);
           M1_WDATABUS         : in   Std_logic_vector(size-1 downto 0);

           -- M2 port
           M2_BUSY,M2_MR,M2_MW : in   Std_logic;
           M2_NREADY           : out  Std_logic;
           M2_ADDRBUS          : in   Std_logic_vector(addr_size-1 downto 0);
           M2_RDATABUS         : out  Std_logic_vector(size-1 downto 0);
           M2_WDATABUS         : in   Std_logic_vector(size-1 downto 0);
		   
           -- S1 port
           S1_BUSY,S1_MR,S1_MW : out  Std_logic;               
           S1_NREADY           : in   Std_logic;
           S1_ADDRBUS          : out  Std_logic_vector(addr_size-1 downto 0);
           S1_RDATABUS         : in   Std_logic_vector(size-1 downto 0);
           S1_WDATABUS         : out  Std_logic_vector(size-1 downto 0);
  
           -- S2 port
           S2_BUSY,S2_MR,S2_MW : out  Std_logic;
           S2_NREADY           : in   Std_logic;
           S2_ADDRBUS          : out  Std_logic_vector(addr_size-1 downto 0);
           S2_RDATABUS         : in   Std_logic_vector(size-1 downto 0);
           S2_WDATABUS         : out  Std_logic_vector(size-1 downto 0);
    
           -- S3 port
           S3_BUSY,S3_MR,S3_MW : out  Std_logic;
           S3_NREADY           : in   Std_logic;
           S3_ADDRBUS          : out  Std_logic_vector(addr_size-1 downto 0);
           S3_RDATABUS         : in   Std_logic_vector(size-1 downto 0);
           S3_WDATABUS         : out  Std_logic_vector(size-1 downto 0);
  
           -- S4 port
           S4_BUSY,S4_MR,S4_MW : out  Std_logic;
           S4_NREADY           : in   Std_logic;
           S4_ADDRBUS          : out  Std_logic_vector(addr_size-1 downto 0);
           S4_RDATABUS         : in   Std_logic_vector(size-1 downto 0);
           S4_WDATABUS         : out  Std_logic_vector(size-1 downto 0) );
  end ubus;

  architecture struct of ubus is

  type master_type is (m1,m2, default);
  type slave_type  is (s1,s2,s3,s4, default);
  type acc_type is (nop, read, write);
      
  type Bus_op is
    record
      master : master_type; 
      slave  : slave_type;
      op     : acc_type;
    end record;

  constant signal_not_active : std_logic := not signal_active;
  signal c1_op,c2_op    : Bus_op;
  signal c1_addrbus     : Std_logic_vector(addr_size-1 downto 0);
  signal c1_nready      : Std_logic;
  signal c1_wdatabus    : Std_logic_vector(size-1 downto 0);
  signal c2_rdatabus    : Std_logic_vector(size-1 downto 0);
  signal c2_busy        : Std_logic;
    
  begin  -- struct

    -- Cycle Bus 1 (Addressing): Determining the prioritary master (priority
    -- policy can be evolved) 
    process(M1_BUSY,M1_MR,M1_MW,M2_BUSY,M2_MR,M2_MW)
    begin
      c1_op.master <= default;
      c1_op.op     <= nop;
      -- Detecting if Master 1 is requiring bus service
      if    (M1_MR=signal_active and M1_BUSY=signal_not_active) then
        c1_op.master <= m1;
        c1_op.op     <= read;
      elsif (M1_MW=signal_active and M1_BUSY=signal_not_active) then
        c1_op.master <= m1;
        c1_op.op     <= write;
      -- Detecting if Master 2 is requiring bus service
      elsif (M2_MR=signal_active and M2_BUSY=signal_not_active) then 
	c1_op.master <= m2;
        c1_op.op     <= read;
      elsif (M2_MW=signal_active and M2_BUSY=signal_not_active) then
        c1_op.master <= m2;
        c1_op.op     <= write;
      end if;
    end process;

      
    addr_Mux: C1_addrbus  <=  M1_ADDRBUS when c1_op.master=m1 else 
                              M2_ADDRBUS when c1_op.master=m2 else 
                              (others=>'0');
				  
    wdata_Mux: C1_wdatabus <= M1_WDATABUS when (c1_op.master=m1 and c1_op.op=write) else 
                              M2_WDATABUS when (c1_op.master=m2 and c1_op.op=write) else
                              (others=>'0');
    
                        
    -- Cycle Bus 1 (Addressing): Determining the Slave to be addressed based on the bus address table
    process(C1_addrbus,c1_op)    
    begin
        c1_op.slave <= default;
        if c1_op.op /= nop then
          if    (unsigned(C1_addrbus) >= resize(unsigned(s1_start),addr_size) ) and
                (unsigned(C1_addrbus) <  resize(unsigned(s1_end),  addr_size) ) then
              c1_op.slave <= s1;          
          elsif (unsigned(C1_addrbus) >= resize(unsigned(s2_start),addr_size) ) and
                (unsigned(C1_addrbus) <  resize(unsigned(s2_end)  ,addr_size) ) then
              c1_op.slave <= s2;       
          elsif (unsigned(C1_addrbus) >= resize(unsigned(s3_start),addr_size)  ) and
                (unsigned(C1_addrbus) <  resize(unsigned(s3_end),  addr_size)  ) then
              c1_op.slave <= s3; 
          elsif (unsigned(C1_addrbus) >= resize(unsigned(s4_start),addr_size) ) and
                (unsigned(C1_addrbus) <  resize(unsigned(s4_end)  ,addr_size) ) then
              c1_op.slave <= s4; 
          end if;
        end if;
    end process;

    -- Still in Cycle Bus 1 (addressing): based on the selected master and the
    -- addressed slave, back-annotation of the appropriate NREADY signal
    c1_nready <=  S1_NREADY when c1_op.slave=s1 else
                  S2_NREADY when c1_op.slave=s2 else
                  S3_NREADY when c1_op.slave=s3 else
                  S4_NREADY when c1_op.slave=s4 else
                 signal_not_active;
    -- NREADY can be asserted in three cases:
    -- a) Master is requiring the bus but another master is having it
    -- b) The slave addressed by the master needs an extension during the addressing
    -- c) The Master in charge of the previous bus run needs an extension during reading
    M1_NREADY   <= signal_active when (M1_MW=signal_active or M1_MR=signal_active) and
                     M1_BUSY=signal_not_active and c1_op.master/=m1 else
                   signal_active when (c1_op.master=m1 and c1_nready=signal_active) else
                   signal_active when (c2_op.master=m2 and M2_BUSY=signal_active) else
                   signal_not_active;
    M2_NREADY   <= signal_active when (M2_MW=signal_active or M2_MR=signal_active) and
                                       M2_BUSY=signal_not_active and c1_op.master/=m2 else
                   signal_active when (c1_op.master=m2 and c1_nready=signal_active) else
                   signal_active when (c2_op.master=m1 and M1_BUSY=signal_active) else                   
                   signal_not_active;
      
    S1_ADDRBUS <= C1_addrbus when c1_op.slave = s1 else (others=>'0');
    S2_ADDRBUS <= C1_addrbus when c1_op.slave = s2 else (others=>'0');
    S3_ADDRBUS <= C1_addrbus when c1_op.slave = s3 else (others=>'0');                   
    S4_ADDRBUS <= C1_addrbus when c1_op.slave = s4 else (others=>'0');

    S1_WDATABUS <= C1_wdatabus when c1_op.slave = s1 else (others=>'0');
    S2_WDATABUS <= C1_wdatabus when c1_op.slave = s2 else (others=>'0');
    S3_WDATABUS <= C1_wdatabus when c1_op.slave = s3 else (others=>'0');
    S4_WDATABUS <= C1_wdatabus when c1_op.slave = s4 else (others=>'0');
    
    S1_MR <= signal_active when c1_op.op=read and c1_op.slave = s1 else signal_not_active;
    S2_MR <= signal_active when c1_op.op=read and c1_op.slave = s2 else signal_not_active;
    S3_MR <= signal_active when c1_op.op=read and c1_op.slave = s3 else signal_not_active;
    S4_MR <= signal_active when c1_op.op=read and c1_op.slave = s4 else signal_not_active;

    S1_MW <= signal_active when c1_op.op=write and c1_op.slave = s1 else signal_not_active;
    S2_MW <= signal_active when c1_op.op=write and c1_op.slave = s2 else signal_not_active;
    S3_MW <= signal_active when c1_op.op=write and c1_op.slave = s3 else signal_not_active;
    S4_MW <= signal_active when c1_op.op=write and c1_op.slave = s4 else signal_not_active;
      
    -- Sequential process sampling the incoming Address in order to route the
    -- relative data upon reading.
    -- Note: here we need to implement eventual waitstates. If the addressed
    -- slave is not ready, we stay in cycle1 and we can't step on to the
    -- following stage. The active master is stalled as well  
    process(clk,reset)
    begin
        if reset='0' then
          C2_op.op <= nop;
          C2_op.master <= default;
          C2_op.slave  <= default;
        else
            if clk'event and clk='1' then
                if c1_nready = signal_not_active then
                    C2_op.op     <= c1_op.op;
                    C2_op.master <= c1_op.master;
                    C2_op.slave  <= c1_op.slave;
                end if;
            end if;
        end if;
    end process;

    -- selecting input value from All slaves
    c2_rdatabus <= S1_RDATABUS when (c2_op.slave=s1 and c2_op.op=read) else
                   S2_RDATABUS when (c2_op.slave=s2 and c2_op.op=read) else
                   S3_RDATABUS when (c2_op.slave=s3 and c2_op.op=read) else
                   S4_RDATABUS when (c2_op.slave=s4 and c2_op.op=read) else
                   (others=> '0');

    c2_busy  <= M1_BUSY when c2_op.master=m1 and c2_op.op=read else
                M2_BUSY when c2_op.master=m2 and c2_op.op=read else
                signal_not_active;   
    
    M1_RDATABUS <= C2_rdatabus when c2_op.master=m1 else (others=>'0');
    M2_RDATABUS <= C2_rdatabus when c2_op.master=m2 else (others=>'0');
  
    S1_BUSY <= c2_busy when c2_op.slave = s1 else signal_not_active;
    S2_BUSY <= c2_busy when c2_op.slave = s2 else signal_not_active;
    S3_BUSY <= c2_busy when c2_op.slave = s3 else signal_not_active;
    S4_BUSY <= c2_busy when c2_op.slave = s4 else signal_not_active;      

  end struct;
